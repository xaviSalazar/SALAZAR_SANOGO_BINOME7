  --Example instantiation for system 'mon_sopc'
  mon_sopc_inst : mon_sopc
    port map(
      AffCentaine_from_the_avalon_gestion_anemo_0 => AffCentaine_from_the_avalon_gestion_anemo_0,
      AffDizane_from_the_avalon_gestion_anemo_0 => AffDizane_from_the_avalon_gestion_anemo_0,
      AffUnite_from_the_avalon_gestion_anemo_0 => AffUnite_from_the_avalon_gestion_anemo_0,
      BCD7SEGMENT_from_the_avalon_gestion_anemo_0 => BCD7SEGMENT_from_the_avalon_gestion_anemo_0,
      data_anemometre_from_the_avalon_gestion_anemo_0 => data_anemometre_from_the_avalon_gestion_anemo_0,
      data_valid_from_the_avalon_gestion_anemo_0 => data_valid_from_the_avalon_gestion_anemo_0,
      done_probe_from_the_avalon_nmea_tx_0 => done_probe_from_the_avalon_nmea_tx_0,
      leds_config_from_the_avalon_gestion_anemo_0 => leds_config_from_the_avalon_gestion_anemo_0,
      multiplex_from_the_avalon_gestion_anemo_0 => multiplex_from_the_avalon_gestion_anemo_0,
      out_pwm_from_the_avalon_pwm_0 => out_pwm_from_the_avalon_pwm_0,
      txd_from_the_avalon_nmea_tx_0 => txd_from_the_avalon_nmea_tx_0,
      val_chaine_from_the_avalon_nmea_rx_0 => val_chaine_from_the_avalon_nmea_rx_0,
      val_data_from_the_avalon_nmea_rx_0 => val_data_from_the_avalon_nmea_rx_0,
      clk_0 => clk_0,
      in_freq_anemometre_to_the_avalon_gestion_anemo_0 => in_freq_anemometre_to_the_avalon_gestion_anemo_0,
      in_port_to_the_switchs_config => in_port_to_the_switchs_config,
      reset_n => reset_n,
      rxd_to_the_avalon_nmea_rx_0 => rxd_to_the_avalon_nmea_rx_0
    );


