  --Example instantiation for system 'mon_sopc'
  mon_sopc_inst : mon_sopc
    port map(
      AffCentaine_from_the_avalon_gestion_anemo_0 => AffCentaine_from_the_avalon_gestion_anemo_0,
      AffDizane_from_the_avalon_gestion_anemo_0 => AffDizane_from_the_avalon_gestion_anemo_0,
      AffUnite_from_the_avalon_gestion_anemo_0 => AffUnite_from_the_avalon_gestion_anemo_0,
      data_anemometre_from_the_avalon_gestion_anemo_0 => data_anemometre_from_the_avalon_gestion_anemo_0,
      data_valid_from_the_avalon_gestion_anemo_0 => data_valid_from_the_avalon_gestion_anemo_0,
      leds_config_from_the_avalon_gestion_anemo_0 => leds_config_from_the_avalon_gestion_anemo_0,
      out_pwm_from_the_avalon_pwm_0 => out_pwm_from_the_avalon_pwm_0,
      clk_0 => clk_0,
      in_freq_anemometre_to_the_avalon_gestion_anemo_0 => in_freq_anemometre_to_the_avalon_gestion_anemo_0,
      in_port_to_the_switchs_config => in_port_to_the_switchs_config,
      reset_n => reset_n
    );


